`timescale 1ns/100ps



module tb

// Uhhhhh mf uhhhh





endmodule