

module matmul #() ();




endmodule




