module tb;





// Test bin2gray function


// Test gray2bin function



endmodule;