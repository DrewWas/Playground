

module tb;

    // Test out multiple dimensions (square, tall, wide etc.)
    // Change N,M,J,K to test non-square matrices


endmodule 