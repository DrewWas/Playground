

module tb;



endmodule 