module tb;





// Test bin2gray function


// Test gray2bin function

// Test at multiple different clks for both read and write 

// Stress test




endmodule;