module and_gate(

    input_1,
    input_2,
    out);


    input input_1;
    input input_2;
    output out;

    assign out = input_1 & input_2;

endmodule

